netcdf cltAnom_rcp85_land-prob_uk_25km_cdf_b8100_1y_mon_19601201-19611130 {
dimensions:
	time = UNLIMITED ; // (12 currently)
	projection_y_coordinate = 52 ;
	projection_x_coordinate = 39 ;
	percentile = 111 ;
	bnds = 2 ;
variables:
	float cltAnom(time, projection_y_coordinate, projection_x_coordinate, percentile) ;
		cltAnom:_FillValue = 1.e+20f ;
		cltAnom:standard_name = "cloud_area_fraction" ;
		cltAnom:long_name = "Cloud area fraction" ;
		cltAnom:units = "%" ;
		cltAnom:anomaly_type = "percentage_change" ;
		cltAnom:description = "Total cloud" ;
		cltAnom:label_units = "%" ;
		cltAnom:plot_label = "Total cloud anomaly (%)" ;
		cltAnom:cell_methods = "time: mean" ;
		cltAnom:grid_mapping = "transverse_mercator" ;
		cltAnom:coordinates = "latitude longitude month_number season_year year" ;
	int transverse_mercator ;
		transverse_mercator:grid_mapping_name = "transverse_mercator" ;
		transverse_mercator:longitude_of_prime_meridian = 0. ;
		transverse_mercator:semi_major_axis = 6377563.396 ;
		transverse_mercator:semi_minor_axis = 6356256.909 ;
		transverse_mercator:longitude_of_central_meridian = -2. ;
		transverse_mercator:latitude_of_projection_origin = 49. ;
		transverse_mercator:false_easting = 400000. ;
		transverse_mercator:false_northing = -100000. ;
		transverse_mercator:scale_factor_at_central_meridian = 0.9996012717 ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:axis = "Y" ;
		projection_y_coordinate:bounds = "projection_y_coordinate_bnds" ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
	double projection_y_coordinate_bnds(projection_y_coordinate, bnds) ;
	int projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:axis = "X" ;
		projection_x_coordinate:bounds = "projection_x_coordinate_bnds" ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
	double projection_x_coordinate_bnds(projection_x_coordinate, bnds) ;
	double percentile(percentile) ;
		percentile:units = "%" ;
		percentile:long_name = "percentile" ;
	double latitude(projection_y_coordinate, projection_x_coordinate) ;
		latitude:units = "1" ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
	double longitude(projection_y_coordinate, projection_x_coordinate) ;
		longitude:units = "1" ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	int season_year(time) ;
		season_year:units = "1" ;
		season_year:long_name = "season_year" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:baseline_period = "b8100" ;
		:collection = "land-prob" ;
		:contact = "ukcpproject@metoffice.gov.uk, UKCP Team, Met Office Hadley Centre" ;
		:creation_date = "2018-10-08T08:34:56" ;
		:domain = "uk" ;
		:frequency = "mon" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:prob_data_type = "cdf" ;
		:project = "UKCP18" ;
		:references = "http://ukclimateprojections.metoffice.gov.uk/" ;
		:resolution = "25km" ;
		:scenario = "rcp85" ;
		:source = "Probabilistic climate prediction based on family of Met Office Hadley Centre climate models HadCM3, HadRM3 and HadSM3, plus climate models from other climate centres contributing to IPCC AR5 and CFMIP." ;
		:time_slice_type = "1y" ;
		:title = "UKCP18 probabilistic projections for total cloud anomaly (%) for UK land points, for the RCP 8.5 scenario with a 1981-2000 baseline." ;
		:version = "v20181004" ;
		:Conventions = "CF-1.5" ;
}
