netcdf psl_rcp85_land-gcm_uk_country_01_ann-30y_196012-199011 {
dimensions:
	ensemble_member = 1 ;
	region = 8 ;
	string24 = 24 ;
	string27 = 27 ;
	bnds = 2 ;
variables:
	float psl(ensemble_member, region) ;
		psl:standard_name = "air_pressure_at_sea_level" ;
		psl:long_name = "Pressure at mean sea level" ;
		psl:units = "hPa" ;
		psl:description = "Sea level pressure" ;
		psl:label_units = "hPa" ;
		psl:plot_label = "Sea level pressure (hPa)" ;
		psl:cell_methods = "time: mean" ;
		psl:coordinates = "ensemble_member_id geo_region time year" ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	char geo_region(region, string24) ;
		geo_region:units = "1" ;
		geo_region:long_name = "Country" ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	double time ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(bnds) ;
	int year ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:collection = "land-gcm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2018-11-22T23:14:33" ;
		:domain = "uk" ;
		:frequency = "ann-30y" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "country" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 global realisation from a set of 15 perturbed variants of HadGEM3-GC3.05 and 13 CMIP5 members that passed a qualitative evaluation" ;
		:title = "UKCP18 land projections - 60km global climate model, sea level pressure (hpa) over the UK for the RCP 8.5 scenario" ;
		:version = "v20181122" ;
		:Conventions = "CF-1.5" ;
}
