netcdf ESACCI-SEAICE-L3C-SITHICK-RA2_ENVISAT-SH50KMEASE2-201202-fv2.0 {
dimensions:
	time = UNLIMITED ; // (1 currently)
	yc = 216 ;
	xc = 216 ;
	nv = 2 ;
variables:
	float freeboard(time, yc, xc) ;
		freeboard:coordinates = "time lon lat" ;
		freeboard:grid_mapping = "Lambert_Azimuthal_Grid" ;
		freeboard:long_name = "elevation of retracked point above instantaneous sea surface height (with snow range corrections)" ;
		freeboard:standard_name = "sea_ice_freeboard" ;
		freeboard:units = "m" ;
	float freeboard_uncertainty(time, yc, xc) ;
		freeboard_uncertainty:coordinates = "time lon lat" ;
		freeboard_uncertainty:grid_mapping = "Lambert_Azimuthal_Grid" ;
		freeboard_uncertainty:long_name = "freeboard uncertainty" ;
		freeboard_uncertainty:units = "m" ;
	double lat(yc, xc) ;
		lat:long_name = "latitude of grid cell center" ;
		lat:standard_name = "latitude" ;
		lat:units = "degrees_north" ;
	double lon(yc, xc) ;
		lon:long_name = "longitude of grid cell center" ;
		lon:standard_name = "longitude" ;
		lon:units = "degrees_east" ;
	float radar_freeboard(time, yc, xc) ;
		radar_freeboard:coordinates = "time lon lat" ;
		radar_freeboard:grid_mapping = "Lambert_Azimuthal_Grid" ;
		radar_freeboard:long_name = "elevation of retracked point above instantaneous sea surface height (no snow range corrections)" ;
		radar_freeboard:units = "m" ;
	float radar_freeboard_uncertainty(time, yc, xc) ;
		radar_freeboard_uncertainty:coordinates = "time lon lat" ;
		radar_freeboard_uncertainty:grid_mapping = "Lambert_Azimuthal_Grid" ;
		radar_freeboard_uncertainty:long_name = "uncertainty of radar freeboard" ;
		radar_freeboard_uncertainty:units = "m" ;
	float sea_ice_concentration(time, yc, xc) ;
		sea_ice_concentration:comment = "Average grid cell sea ice concentration during days with altimetry data coverage (not monthly mean)" ;
		sea_ice_concentration:coordinates = "time lon lat" ;
		sea_ice_concentration:grid_mapping = "Lambert_Azimuthal_Grid" ;
		sea_ice_concentration:long_name = "sea ice contration" ;
		sea_ice_concentration:standard_name = "sea_ice_area_fraction" ;
		sea_ice_concentration:units = "percent" ;
		sea_ice_concentration:valid_max = 100. ;
		sea_ice_concentration:valid_min = 0. ;
	float sea_ice_thickness(time, yc, xc) ;
		sea_ice_thickness:ancillary_variables = "sea_ice_thickness_uncertainty status_flag" ;
		sea_ice_thickness:coordinates = "time lon lat" ;
		sea_ice_thickness:grid_mapping = "Lambert_Azimuthal_Grid" ;
		sea_ice_thickness:long_name = "thickness of the sea ice layer" ;
		sea_ice_thickness:standard_name = "sea_ice_thickness" ;
		sea_ice_thickness:units = "m" ;
	float sea_ice_thickness_uncertainty(time, yc, xc) ;
		sea_ice_thickness_uncertainty:coordinates = "time lon lat" ;
		sea_ice_thickness_uncertainty:grid_mapping = "Lambert_Azimuthal_Grid" ;
		sea_ice_thickness_uncertainty:long_name = "uncertainty of the sea ice layer thickness" ;
		sea_ice_thickness_uncertainty:units = "m" ;
	byte status_flag(time, yc, xc) ;
		status_flag:comment = "Describes the status of the sea-ice thickness retrieval" ;
		status_flag:coordinates = "time lat lon" ;
		status_flag:flag_meaning = "0: nominal sea ice thickness retrieval; 1: no input data; 2: outside sea ice concentration mask; 3: latitude above orbit inclination; 4: land, lake or land ice; 5: sea ice thickness retrieval failed;" ;
		status_flag:flag_values = 0, 1, 2, 3, 4, 5 ;
		status_flag:grid_mapping = "Lambert_Azimuthal_Grid" ;
		status_flag:long_name = "status flag for the sea ice thickness retrieval" ;
		status_flag:standard_name = "sea_ice_thickness status_flag" ;
		status_flag:unit = 1 ;
		status_flag:valid_max = 5 ;
		status_flag:valid_min = 0 ;
	double time(time) ;
		time:standard_name = "time" ;
		time:units = "seconds since 1970-01-01" ;
		time:long_name = "reference time of product" ;
		time:axis = "T" ;
		time:calendar = "standard" ;
		time:bounds = "time_bnds" ;
	double time_bnds(time, nv) ;
		time_bnds:units = "seconds since 1970-01-01" ;
	double xc(xc) ;
		xc:standard_name = "projection_x_coordinate" ;
		xc:units = "km" ;
		xc:long_name = "x coordinate of projection (eastings)" ;
	double yc(yc) ;
		yc:standard_name = "projection_y_coordinate" ;
		yc:units = "km" ;
		yc:long_name = "y coordinate of projection (eastings)" ;
	byte Lambert_Azimuthal_Grid ;
		Lambert_Azimuthal_Grid:false_easting = 0. ;
		Lambert_Azimuthal_Grid:false_northing = 0. ;
		Lambert_Azimuthal_Grid:grid_mapping_name = "lambert_azimuthal_equal_area" ;
		Lambert_Azimuthal_Grid:inverse_flattening = 298.257223563 ;
		Lambert_Azimuthal_Grid:latitude_of_projection_origin = -90. ;
		Lambert_Azimuthal_Grid:longitude_of_projection_origin = 0. ;
		Lambert_Azimuthal_Grid:proj4_string = "+proj=laea +lon_0=0 +datum=WGS84 +ellps=WGS84 +lat_0=-90.0" ;
		Lambert_Azimuthal_Grid:semi_major_axis = 6378137. ;

// global attributes:
		:title = "ESA Climate Change Initiative Sea Ice: Experimental Southern Hemisphere Sea Ice Thickness Climate Data Record" ;
		:institution = "Alfred-Wegener-Institut Helmholtz Zentrum für Polar und Meeresforschung" ;
		:source = "Altimetry: envisat, Snow depth: ESA-SICCI AMSR-E/AMSR2 snow depth on sea ice climatology, Mean Sea Surface: DTU15 global mean sea surface, Sea ice Concentration: OSI-SAF Global Sea Ice Concentration (OSI-409), Sea ice type:  First-year sea ice only" ;
		:platform = "Envisat" ;
		:sensor = "RA-2" ;
		:history = "20180417T184311Z (created)" ;
		:references = "Algorithm Theoretical Baseline Document, Sea Ice Climate Change Initiative: Phase 2 (version 2.2)" ;
		:tracking_id = "1a6cb716-a7ba-4c8b-89a3-b601c96520e1" ;
		:conventions = "CF-1.6" ;
		:product_version = "2.0" ;
		:processing_level = "Level-3 Collated (l3c)" ;
		:summary = "Monthly gridded Southern Hemisphere Sea Ice Thickness Climate Data Record from Envisat and CryoSat-2 satellite radar altimetry for the period June 2002 - April 2017." ;
		:keywords = "Sea Ice, Ice Depth/Thickness, Radar Altimeters" ;
		:id = "esacci-seaice-l3c-sit-RA-2-envisat-sh50kmEASE2-20120201-fv2.0" ;
		:naming_authority = "de.awi" ;
		:keywords_vocabulary = "GCMD Science Keywords" ;
		:doi = "10.5285/b1f1ac03077b4aa784c5a413a2210bf5" ;
		:cdm_data_type = "Grid" ;
		:comment = "Southern hemisphere sea ice thickness is an experimental climate data record, as the algorithm does not properly considers the impact of the complex snow morphology in the freeboard retrieval. Sea ice thickness is provided for all month but needs to be considered biased high in areas with high snow depth and during the southern summer month. Please consult the Product User Guide (PUG) for more information." ;
		:date_created = "20180417T184311Z" ;
		:creator_name = "Stefan Hendricks, Stephan Paul (Alfred Wegener Institute Helmholtz Centre for Polar and Marine Research, Bremerhaven, Germany); Eero Rine (Finnish Meteorological Institute, Helsinki, Finland)" ;
		:creator_url = "http://www.awi.de" ;
		:creator_email = "stefan.hendricks@awi.de, stephan.paul@awi.de, eero.rinne@fmi.fi" ;
		:project = "Climate Change Initiative - European Space Agency" ;
		:geospatial_lat_min = "-89.6835" ;
		:geospatial_lat_max = "-16.8229" ;
		:geospatial_lon_min = "-179.7335" ;
		:geospatial_lon_max = "179.7335" ;
		:geospatial_vertical_min = "0.0" ;
		:geospatial_vertical_max = "0.0" ;
		:time_coverage_start = "20120201T000000Z" ;
		:time_coverage_end = "20120229T235959Z" ;
		:time_coverage_duration = "P1M" ;
		:time_coverage_resolution = "P1M" ;
		:spatial_resolution = "50 km" ;
		:standard_name_vocabulary = "CF" ;
		:license = "Creative Commons Attribution 4.0 International (CC BY 4.0)" ;
}
