netcdf pslAnom_rcp85_land-prob_uk_river_pdf_b8110_30y_mon_20091201-20991130 {
dimensions:
	time = 84 ;
	region = 23 ;
	percentile = 111 ;
	bnds = 2 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float pslAnom(time, region, percentile) ;
		pslAnom:long_name = "Pressure at mean sea level" ;
		pslAnom:units = "hPa" ;
		pslAnom:anomaly_type = "absolute_change" ;
		pslAnom:description = "Sea level pressure" ;
		pslAnom:label_units = "hPa-1" ;
		pslAnom:plot_label = "Probability density for sea level pressure anomaly (hPa-1)" ;
		pslAnom:cell_methods = "time: mean" ;
		pslAnom:coordinates = "geo_region month_number season season_year year" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	double percentile(percentile) ;
		percentile:units = "%" ;
		percentile:long_name = "percentile" ;
	char geo_region(region, string27) ;
		geo_region:units = "no_unit" ;
		geo_region:long_name = "River Basin" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	char season(time, string64) ;
		season:units = "1" ;
		season:long_name = "season" ;
	int season_year(time) ;
		season_year:units = "1" ;
		season_year:long_name = "season_year" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:baseline_period = "b8110" ;
		:collection = "land-prob" ;
		:contact = "ukcpproject@metoffice.gov.uk, UKCP Team, Met Office Hadley Centre" ;
		:creation_date = "2018-12-23T16:07:17" ;
		:domain = "uk" ;
		:frequency = "mon" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:prob_data_type = "pdf" ;
		:project = "UKCP18" ;
		:references = "http://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "river" ;
		:scenario = "rcp85" ;
		:source = "Probabilistic climate prediction based on family of Met Office Hadley Centre climate models HadCM3, HadRM3 and HadSM3, plus climate models from other climate centres contributing to IPCC AR5 and CFMIP." ;
		:time_slice_type = "30y" ;
		:title = "UKCP18 probabilistic projections for sea level pressure anomaly (hPa) for UK land points, for the RCP 8.5 scenario with a 1981-2010 baseline." ;
		:version = "v20181122" ;
		:Conventions = "CF-1.5" ;
}
