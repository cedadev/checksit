netcdf tasmax_rcp85_land-rcm_uk_12km_EC-EARTH_r12i1p1_HIRHAM5_day_19801201-19901130 {
dimensions:
	ensemble_member = 1 ;
	projection_y_coordinate = 112 ;
	projection_x_coordinate = 82 ;
	time = 3652 ;
	bnds = 2 ;
	string46 = 46 ;
	string64 = 64 ;
variables:
	string ensemble_member(ensemble_member) ;
	double projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:_FillValue = NaN ;
		projection_y_coordinate:axis = "Y" ;
		projection_y_coordinate:bounds = "projection_y_coordinate_bnds" ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
	double projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:_FillValue = NaN ;
		projection_x_coordinate:axis = "X" ;
		projection_x_coordinate:bounds = "projection_x_coordinate_bnds" ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
	double time(time) ;
		time:_FillValue = NaN ;
		time:standard_name = "time" ;
		time:bounds = "time_bnds" ;
		time:long_name = "time" ;
		time:cell_methods = "time: mean" ;
		time:units = "days since 1949-12-01" ;
		time:calendar = "proleptic_gregorian" ;
	double tasmax(ensemble_member, time, projection_y_coordinate, projection_x_coordinate) ;
		tasmax:_FillValue = NaN ;
		tasmax:regrid_method = "conservative_normed" ;
		tasmax:grid_mapping = "transverse_mercator" ;
		tasmax:coordinates = "grid_longitude month_number grid_latitude ensemble_member_id year yyyymmdd" ;
	int transverse_mercator ;
		transverse_mercator:grid_mapping_name = "transverse_mercator" ;
		transverse_mercator:longitude_of_prime_meridian = 0. ;
		transverse_mercator:semi_major_axis = 6377563.396 ;
		transverse_mercator:semi_minor_axis = 6356256.909 ;
		transverse_mercator:longitude_of_central_meridian = -2. ;
		transverse_mercator:latitude_of_projection_origin = 49. ;
		transverse_mercator:false_easting = 400000. ;
		transverse_mercator:false_northing = -100000. ;
		transverse_mercator:scale_factor_at_central_meridian = 0.9996012717 ;
	int64 time_bnds(time, bnds) ;
		time_bnds:coordinates = "year yyyymmdd month_number" ;
	double projection_y_coordinate_bnds(projection_y_coordinate, bnds) ;
		projection_y_coordinate_bnds:_FillValue = NaN ;
	double projection_x_coordinate_bnds(projection_x_coordinate, bnds) ;
		projection_x_coordinate_bnds:_FillValue = NaN ;
	char ensemble_member_id(ensemble_member, string46) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	double grid_longitude(projection_y_coordinate, projection_x_coordinate) ;
		grid_longitude:_FillValue = NaN ;
		grid_longitude:units = "degrees_east" ;
		grid_longitude:standard_name = "grid_longitude" ;
	double grid_latitude(projection_y_coordinate, projection_x_coordinate) ;
		grid_latitude:_FillValue = NaN ;
		grid_latitude:units = "degrees_north" ;
		grid_latitude:standard_name = "grid_latitude" ;
	int64 month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	int64 year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;
	char yyyymmdd(time, string64) ;
		yyyymmdd:units = "1" ;
		yyyymmdd:long_name = "yyyymmdd" ;

// global attributes:
		:collection = "EuroCORDEX" ;
		:contact = "clair.barnes.16@ucl.ac.uk" ;
		:creation_date = "2022-02-08T16:25:09" ;
		:domain = "uk" ;
		:frequency = "day" ;
		:institution = "Danish Meteorological Institute" ;
		:institution_id = "DMI" ;
		:project = "CORDEX" ;
		:resolution = "12km" ;
		:scenario = "rcp85" ;
		:source = "EuroCORDEX downscaled climate projections based on historical + rcp85 scenarios." ;
		string :title = "EuroCORDEX regional projections for maximum air temperature at 1.5m (°C) for the UK, for the historical + RCP 8.5 scenarios." ;
		:version = "" ;
		:Conventions = "CF-1.6" ;
		:driving_model_id = "ICHEC-EC-EARTH" ;
		:model_id = "DMI-HIRHAM5" ;
		:driving_model_ensemble_member = "r12i1p1" ;
		:rcm_version_id = "v1" ;
}
