netcdf clt_rcp85_land-gcm_uk_country_01_mon_189912-209911 {
dimensions:
	ensemble_member = 1 ;
	time = 2400 ;
	region = 8 ;
	bnds = 2 ;
	string24 = 24 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float clt(ensemble_member, time, region) ;
		clt:standard_name = "cloud_area_fraction" ;
		clt:long_name = "Cloud area fraction" ;
		clt:units = "%" ;
		clt:description = "Total cloud" ;
		clt:label_units = "%" ;
		clt:plot_label = "Total cloud (%)" ;
		clt:cell_methods = "time: mean" ;
		clt:coordinates = "ensemble_member_id geo_region month_number year yyyymm" ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	char geo_region(region, string24) ;
		geo_region:units = "1" ;
		geo_region:long_name = "Country" ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;
	char yyyymm(time, string64) ;
		yyyymm:units = "1" ;
		yyyymm:long_name = "yyyymm" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:collection = "land-gcm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2018-11-05T13:58:58" ;
		:domain = "uk" ;
		:frequency = "mon" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "country" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 global realisation from a set of 15 perturbed variants of HadGEM3-GC3.05 and 13 CMIP5 members that passed a qualitative evaluation" ;
		:title = "UKCP18 land projections - 60km global climate model, total cloud (%) over the UK for the RCP 8.5 scenario" ;
		:version = "v20181122" ;
		:Conventions = "CF-1.5" ;
}
