netcdf uas_rcp85_land-rcm_uk_12km_01_ann-20y_198012-200011 {
dimensions:
	ensemble_member = 1 ;
	projection_y_coordinate = 112 ;
	projection_x_coordinate = 82 ;
	bnds = 2 ;
	string27 = 27 ;
variables:
	float uas(ensemble_member, projection_y_coordinate, projection_x_coordinate) ;
		uas:_FillValue = 1.e+20f ;
		uas:standard_name = "eastward_wind" ;
		uas:long_name = "Eastward wind component" ;
		uas:units = "m s-1" ;
		uas:description = "Eastward wind" ;
		uas:label_units = "m s-1" ;
		uas:plot_label = "Eastward wind at 10m (m s-1)" ;
		uas:cell_methods = "time: mean" ;
		uas:grid_mapping = "transverse_mercator" ;
		uas:coordinates = "ensemble_member_id grid_latitude grid_longitude time year" ;
	int transverse_mercator ;
		transverse_mercator:grid_mapping_name = "transverse_mercator" ;
		transverse_mercator:longitude_of_prime_meridian = 0. ;
		transverse_mercator:semi_major_axis = 6377563.396 ;
		transverse_mercator:semi_minor_axis = 6356256.909 ;
		transverse_mercator:longitude_of_central_meridian = -2. ;
		transverse_mercator:latitude_of_projection_origin = 49. ;
		transverse_mercator:false_easting = 400000. ;
		transverse_mercator:false_northing = -100000. ;
		transverse_mercator:scale_factor_at_central_meridian = 0.9996012717 ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:axis = "Y" ;
		projection_y_coordinate:bounds = "projection_y_coordinate_bnds" ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
	double projection_y_coordinate_bnds(projection_y_coordinate, bnds) ;
	double projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:axis = "X" ;
		projection_x_coordinate:bounds = "projection_x_coordinate_bnds" ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
	double projection_x_coordinate_bnds(projection_x_coordinate, bnds) ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	double grid_latitude(projection_y_coordinate, projection_x_coordinate) ;
		grid_latitude:units = "degrees_north" ;
		grid_latitude:standard_name = "grid_latitude" ;
	double grid_longitude(projection_y_coordinate, projection_x_coordinate) ;
		grid_longitude:units = "degrees_east" ;
		grid_longitude:standard_name = "grid_longitude" ;
	double time ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(bnds) ;
	int year ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:collection = "land-rcm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2019-07-31T00:00:00" ;
		:domain = "uk" ;
		:frequency = "ann-20y" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "12km" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 regional realisation from a set of 12 limited-area Met Office Unified Model Global Atmosphere GA7 models at 12km resolution driven by perturbed variants of the global HadGEM3-GC3.05" ;
		:title = "UKCP18 land projections - 12km regional climate model, eastward wind at 10m (m s-1) over the UK for the RCP 8.5 scenario" ;
		:version = "v20190731" ;
		:Conventions = "CF-1.5" ;
}
