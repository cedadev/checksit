netcdf rls_rcp85_land-rcm_uk_region_01_ann-30y_198012-201011 {
dimensions:
	ensemble_member = 1 ;
	region = 16 ;
	string24 = 24 ;
	string27 = 27 ;
	bnds = 2 ;
variables:
	float rls(ensemble_member, region) ;
		rls:standard_name = "surface_net_downward_longwave_flux" ;
		rls:long_name = "Net Surface long wave flux" ;
		rls:units = "W m-2" ;
		rls:description = "Net Surface long wave flux" ;
		rls:label_units = "W m-2" ;
		rls:plot_label = "Net Surface long wave flux (W m-2)" ;
		rls:cell_methods = "time: mean" ;
		rls:coordinates = "ensemble_member_id geo_region time year" ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	char geo_region(region, string24) ;
		geo_region:units = "1" ;
		geo_region:long_name = "Region" ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	double time ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(bnds) ;
	int year ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:collection = "land-rcm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2018-11-22T23:15:07" ;
		:domain = "uk" ;
		:frequency = "ann-30y" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "region" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 regional realisation from a set of 12 limited-area Met Office Unified Model Global Atmosphere GA7 models at 12km resolution driven by perturbed variants of the global HadGEM3-GC3.05" ;
		:title = "UKCP18 land projections - 12km regional climate model, net surface long wave flux (w m-2) over the UK for the RCP 8.5 scenario" ;
		:version = "v20181122" ;
		:Conventions = "CF-1.5" ;
}
