netcdf tasmin_rcp85_land-rcm_uk_river_01_day_19801201-20801130 {
dimensions:
	ensemble_member = 1 ;
	time = 36000 ;
	region = 23 ;
	bnds = 2 ;
	string24 = 24 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float tasmin(ensemble_member, time, region) ;
		tasmin:standard_name = "air_temperature" ;
		tasmin:long_name = "Minimum air temperature" ;
		tasmin:units = "degC" ;
		tasmin:description = "Minimum air temperature" ;
		tasmin:label_units = "°C" ;
		tasmin:plot_label = "Minimum air temperature at 1.5m (°C)" ;
		tasmin:cell_methods = "time: minimum" ;
		tasmin:coordinates = "ensemble_member_id geo_region month_number year yyyymmdd" ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	char geo_region(region, string24) ;
		geo_region:units = "1" ;
		geo_region:long_name = "River" ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;
	char yyyymmdd(time, string64) ;
		yyyymmdd:units = "1" ;
		yyyymmdd:long_name = "yyyymmdd" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:collection = "land-rcm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2018-11-10T16:13:28" ;
		:domain = "uk" ;
		:frequency = "day" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "river" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 regional realisation from a set of 12 limited-area Met Office Unified Model Global Atmosphere GA7 models at 12km resolution driven by perturbed variants of the global HadGEM3-GC3.05" ;
		:title = "UKCP18 land projections - 12km regional climate model, minimum air temperature at 1.5m (°c) over the UK for the RCP 8.5 scenario" ;
		:version = "v20181122" ;
		:Conventions = "CF-1.5" ;
}
