netcdf ncas-dewpoint-hygrometer-1_mobile_18600101_dew-point_v1.0 {
dimensions:
	latitude = 1 ;
	longitude = 1 ;
	time = 10 ;
variables:
	float dew_point_temperature(time) ;
		dew_point_temperature:_FillValue = -1.e+20f ;
		dew_point_temperature:units = "K" ;
		dew_point_temperature:standard_name = "dew_point_temperature" ;
		dew_point_temperature:long_name = "Dew \\Frost point Temperature" ;
		dew_point_temperature:valid_min = "<derived from file>" ;
		dew_point_temperature:valid_max = "<derived from file>" ;
		dew_point_temperature:cell_methods = "EXAMPLE: time: mean or time: point" ;
		dew_point_temperature:coordinates = "latitude longitude" ;
	float relative_humidity(time) ;
		relative_humidity:_FillValue = -1.e+20f ;
		relative_humidity:units = "%" ;
		relative_humidity:standard_name = "relative_humidity" ;
		relative_humidity:long_name = "Relative Humidity" ;
		relative_humidity:valid_min = "<derived from file>" ;
		relative_humidity:valid_max = "<derived from file>" ;
		relative_humidity:cell_methods = "EXAMPLE: time: mean or time: point" ;
		relative_humidity:coordinates = "latitude longitude" ;
	float mole_fraction_of_water_vapor_in_air(time) ;
		mole_fraction_of_water_vapor_in_air:_FillValue = -1.e+20f ;
		mole_fraction_of_water_vapor_in_air:units = "EXAMPLE: 1|1e-3|1e-6|1e-9|1e-12" ;
		mole_fraction_of_water_vapor_in_air:practical_units = "EXAMPLE: mmol mol-1|micro mol mol-1|nmol mol-1|pmol mol-1" ;
		mole_fraction_of_water_vapor_in_air:standard_name = "mole_fraction_of_water_vapor_in_air" ;
		mole_fraction_of_water_vapor_in_air:long_name = "Mole Fraction of Water Vapour in air" ;
		mole_fraction_of_water_vapor_in_air:valid_min = "<derived from file>" ;
		mole_fraction_of_water_vapor_in_air:valid_max = "<derived from file>" ;
		mole_fraction_of_water_vapor_in_air:cell_methods = "EXAMPLE: time: mean or time: point" ;
		mole_fraction_of_water_vapor_in_air:coordinates = "latitude longitude" ;
		mole_fraction_of_water_vapor_in_air:chemical_species = "H2O" ;
	float mass_fraction_of_water_vapor_in_air(time) ;
		mass_fraction_of_water_vapor_in_air:_FillValue = -1.e+20f ;
		mass_fraction_of_water_vapor_in_air:units = "EXAMPLE: 1|1e-3|1e-6|1e-9|1e-12" ;
		mass_fraction_of_water_vapor_in_air:practical_units = "EXAMPLE: ppm|ppb|ppt" ;
		mass_fraction_of_water_vapor_in_air:long_name = "Mass Fraction of Water Vapour in air" ;
		mass_fraction_of_water_vapor_in_air:valid_min = "<derived from file>" ;
		mass_fraction_of_water_vapor_in_air:valid_max = "<derived from file>" ;
		mass_fraction_of_water_vapor_in_air:cell_methods = "EXAMPLE: time: mean or time: point" ;
		mass_fraction_of_water_vapor_in_air:coordinates = "latitude longitude" ;
		mass_fraction_of_water_vapor_in_air:chemical_species = "H2O" ;
	float mole_concentration_of_water_vapor_in_air(time) ;
		mole_concentration_of_water_vapor_in_air:_FillValue = -1.e+20f ;
		mole_concentration_of_water_vapor_in_air:units = "mol m-3" ;
		mole_concentration_of_water_vapor_in_air:standard_name = "mole_concentration_of_water_vapor_in_air" ;
		mole_concentration_of_water_vapor_in_air:long_name = "Mole Concentration of Water Vapour in air" ;
		mole_concentration_of_water_vapor_in_air:valid_min = "<derived from file>" ;
		mole_concentration_of_water_vapor_in_air:valid_max = "<derived from file>" ;
		mole_concentration_of_water_vapor_in_air:cell_methods = "EXAMPLE: time: mean or time: point" ;
		mole_concentration_of_water_vapor_in_air:coordinates = "latitude longitude" ;
		mole_concentration_of_water_vapor_in_air:chemical_species = "H2O" ;
	float mass_concentration_of_water_vapor_in_air(time) ;
		mass_concentration_of_water_vapor_in_air:_FillValue = -1.e+20f ;
		mass_concentration_of_water_vapor_in_air:units = "kg m-3" ;
		mass_concentration_of_water_vapor_in_air:standard_name = "mass_concentration_of_water_vapor_in_air" ;
		mass_concentration_of_water_vapor_in_air:long_name = "Mass Concentration of Water Vapour in air" ;
		mass_concentration_of_water_vapor_in_air:valid_min = "<derived from file>" ;
		mass_concentration_of_water_vapor_in_air:valid_max = "<derived from file>" ;
		mass_concentration_of_water_vapor_in_air:cell_methods = "EXAMPLE: time: mean or time: point" ;
		mass_concentration_of_water_vapor_in_air:coordinates = "latitude longitude" ;
		mass_concentration_of_water_vapor_in_air:chemical_species = "H2O" ;
	byte qc_flag(time) ;
		qc_flag:units = "1" ;
		qc_flag:long_name = "Data Quality flag" ;
		qc_flag:flag_values = 0b, 1b, 2b, 3b ;
		qc_flag:flag_meanings = "not_used good_data suspect_data_contact_creator bad_data_do_not_use" ;
	double time(time) ;
		time:units = "seconds since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:long_name = "Time (seconds since 1970-01-01 00:00:00)" ;
		time:axis = "T" ;
		time:valid_min = "<derived from file>" ;
		time:valid_max = "<derived from file>" ;
		time:calendar = "standard" ;
	float latitude(latitude) ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "Latitude" ;
	float longitude(longitude) ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "Longitude" ;
	float day_of_year(time) ;
		day_of_year:units = "1" ;
		day_of_year:long_name = "Day of Year" ;
		day_of_year:valid_min = "<derived from file>" ;
		day_of_year:valid_max = "<derived from file>" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "Year" ;
		year:valid_min = "<derived from file>" ;
		year:valid_max = "<derived from file>" ;
	int month(time) ;
		month:units = "1" ;
		month:long_name = "Month" ;
		month:valid_min = "<derived from file>" ;
		month:valid_max = "<derived from file>" ;
	int day(time) ;
		day:units = "1" ;
		day:long_name = "Day" ;
		day:valid_min = "<derived from file>" ;
		day:valid_max = "<derived from file>" ;
	int hour(time) ;
		hour:units = "1" ;
		hour:long_name = "Hour" ;
		hour:valid_min = "<derived from file>" ;
		hour:valid_max = "<derived from file>" ;
	int minute(time) ;
		minute:units = "1" ;
		minute:long_name = "Minute" ;
		minute:valid_min = "<derived from file>" ;
		minute:valid_max = "<derived from file>" ;
	float second(time) ;
		second:units = "1" ;
		second:long_name = "Second" ;
		second:valid_min = "<derived from file>" ;
		second:valid_max = "<derived from file>" ;

// global attributes:
		:Conventions = "CF-1.6, NCAS-AMF-2.0.0" ;
		:source = "NCAS Dewpoint Hygrometer unit 1" ;
		:instrument_manufacturer = "General Eastern" ;
		:instrument_model = "Optica Chilled Mirror Hygrometer" ;
		:instrument_serial_number = "" ;
		:institution = "National Centre for Atmospheric Science (NCAS)" ;
		:last_revised_date = "2023-08-25T09:01:16" ;
		:licence = "Data usage licence - UK Government Open Licence agreement: http://www.nationalarchives.gov.uk/doc/open-government-licence" ;
		:acknowledgement = "Acknowledgement of NCAS as the data provider is required whenever and wherever these data are used" ;
		:platform = "mobile" ;
		:deployment_mode = "land" ;
		:amf_vocabularies_release = "https://github.com/ncasuk/AMF_CVs/releases/tag/v2.0.0" ;
		:history = "2023-08-25T09:01:16 - File created by earjham on ncas-obs-sci-m-202205131617.ncas-obs-sci-m.jasmin.ac.uk using the ncas_amof_netcdf_template python package" ;
		:comment = "CHANGE: Any other text that might be useful. Use \"None\" if no comment needed.. String: min 4 characters" ;
		:instrument_software = "Instrument software" ;
		:instrument_software_version = "v1" ;
		:creator_name = "Rudolf Clausius" ;
		:creator_email = "rudolf.clausius@ncas.ac.uk" ;
		:creator_url = "n/a" ;
		:processing_software_url = "https://not.github.com/rudolf-clausius/instrument-processing-software" ;
		:processing_software_version = "v1" ;
		:calibration_sensitivity = "close enough" ;
		:calibration_certification_date = "n/a" ;
		:calibration_certification_url = "n/a" ;
		:sampling_interval = "5 seconds" ;
		:averaging_interval = "5 seconds" ;
		:product_version = "v1.0" ;
		:processing_level = 0 ;
		:project = "Historic measurements" ;
		:project_principal_investigator = "Benoit Paul Emile Clapyron" ;
		:project_principal_investigator_email = "emile.clapyron@ncas.ac.uk" ;
		:project_principal_investigator_url = "n/a" ;
		:platform_type = "cao" ;
		:title = "Historic measurements of humidity" ;
		:featureType = "timeSeries" ;
		:time_coverage_start = "1860-01-01T00:00:00" ;
		:time_coverage_end = "1860-01-01T23:59:59" ;
		:geospatial_bounds = "47.376 8.548" ;
		:platform_altitude = "408 m" ;
		:location_keywords = "Zurich" ;
}
