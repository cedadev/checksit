netcdf rss_rcp85_land-cpm_uk_5km_01_day_19801201-19901130 {
dimensions:
	ensemble_member = 1 ;
	time = 3600 ;
	projection_y_coordinate = 244 ;
	projection_x_coordinate = 180 ;
	bnds = 2 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float rss(ensemble_member, time, projection_y_coordinate, projection_x_coordinate) ;
		rss:_FillValue = 1.e+20f ;
		rss:standard_name = "surface_net_downward_shortwave_flux" ;
		rss:long_name = "Net Surface short wave flux" ;
		rss:units = "W m-2" ;
		rss:description = "Net Surface short wave flux" ;
		rss:label_units = "W m-2" ;
		rss:plot_label = "Net Surface short wave flux (W m-2)" ;
		rss:cell_methods = "time: mean" ;
		rss:grid_mapping = "transverse_mercator" ;
		rss:coordinates = "ensemble_member_id latitude longitude month_number year yyyymmdd" ;
	int transverse_mercator ;
		transverse_mercator:grid_mapping_name = "transverse_mercator" ;
		transverse_mercator:longitude_of_prime_meridian = 0. ;
		transverse_mercator:semi_major_axis = 6377563.396 ;
		transverse_mercator:semi_minor_axis = 6356256.909 ;
		transverse_mercator:longitude_of_central_meridian = -2. ;
		transverse_mercator:latitude_of_projection_origin = 49. ;
		transverse_mercator:false_easting = 400000. ;
		transverse_mercator:false_northing = -100000. ;
		transverse_mercator:scale_factor_at_central_meridian = 0.9996012717 ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	double projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:axis = "Y" ;
		projection_y_coordinate:bounds = "projection_y_coordinate_bnds" ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
	double projection_y_coordinate_bnds(projection_y_coordinate, bnds) ;
	double projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:axis = "X" ;
		projection_x_coordinate:bounds = "projection_x_coordinate_bnds" ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
	double projection_x_coordinate_bnds(projection_x_coordinate, bnds) ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	double latitude(projection_y_coordinate, projection_x_coordinate) ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	double longitude(projection_y_coordinate, projection_x_coordinate) ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;
	char yyyymmdd(time, string64) ;
		yyyymmdd:units = "1" ;
		yyyymmdd:long_name = "yyyymmdd" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.6.1|hdf5libversion=1.10.4" ;
		:collection = "land-cpm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2021-06-09T16:58:01" ;
		:domain = "uk" ;
		:frequency = "day" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "5km" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 realisation from a set of 12 convection-permitting models (HadREM3-RA11M) driven by perturbed variants of the Met Office Unified Model Global Atmosphere GA7 model (HadREM3-GA705) at 12km resolution.  The HadREM3-GA705 models were driven by perturbed variants of the global HadGEM3-GC3.05" ;
		:title = "UKCP18 land projections - Regridded 2.2km convection-permitting climate model results on 5km British National Grid from Ordnance Survey (OSGB), Net Surface short wave flux over the UK for the RCP8.5 scenario" ;
		:version = "v20210615" ;
		:Conventions = "CF-1.7" ;
}
