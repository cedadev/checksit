netcdf tasmax_rcp85_land-gcm_uk_region_01_seas-30y_196012-199011 {
dimensions:
	ensemble_member = 1 ;
	time = 4 ;
	region = 16 ;
	bnds = 2 ;
	string24 = 24 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float tasmax(ensemble_member, time, region) ;
		tasmax:standard_name = "air_temperature" ;
		tasmax:long_name = "Maximum air temperature" ;
		tasmax:units = "degC" ;
		tasmax:description = "Maximum air temperature" ;
		tasmax:label_units = "°C" ;
		tasmax:plot_label = "Maximum air temperature at 1.5m (°C)" ;
		tasmax:cell_methods = "time: maximum" ;
		tasmax:coordinates = "ensemble_member_id geo_region season year" ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	char geo_region(region, string24) ;
		geo_region:units = "1" ;
		geo_region:long_name = "Region" ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	char season(time, string64) ;
		season:units = "1" ;
		season:long_name = "season" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:collection = "land-gcm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2018-11-22T23:14:33" ;
		:domain = "uk" ;
		:frequency = "seas-30y" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "region" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 global realisation from a set of 15 perturbed variants of HadGEM3-GC3.05 and 13 CMIP5 members that passed a qualitative evaluation" ;
		:title = "UKCP18 land projections - 60km global climate model, maximum air temperature at 1.5m (°c) over the UK for the RCP 8.5 scenario" ;
		:version = "v20181122" ;
		:Conventions = "CF-1.5" ;
}
