netcdf hussAnom_rcp85_land-prob_uk_river_cdf_b8100_1y_mon_19601201-20991130 {
dimensions:
	time = UNLIMITED ; // (1668 currently)
	region = 23 ;
	percentile = 111 ;
	bnds = 2 ;
	string27 = 27 ;
variables:
	float hussAnom(time, region, percentile) ;
		hussAnom:standard_name = "specific_humidity" ;
		hussAnom:long_name = "Specific humidity" ;
		hussAnom:units = "%" ;
		hussAnom:anomaly_type = "percentage_change" ;
		hussAnom:description = "Specific humidity" ;
		hussAnom:label_units = "%" ;
		hussAnom:plot_label = "Specific humidity anomaly at 1.5m (%)" ;
		hussAnom:cell_methods = "time: mean" ;
		hussAnom:coordinates = "geo_region month_number year" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	double percentile(percentile) ;
		percentile:units = "%" ;
		percentile:long_name = "percentile" ;
	char geo_region(region, string27) ;
		geo_region:units = "1" ;
		geo_region:long_name = "River Basin" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:baseline_period = "b8100" ;
		:collection = "land-prob" ;
		:contact = "ukcpproject@metoffice.gov.uk, UKCP Team, Met Office Hadley Centre" ;
		:creation_date = "2018-12-23T16:07:17" ;
		:domain = "uk" ;
		:frequency = "mon" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:prob_data_type = "cdf" ;
		:project = "UKCP18" ;
		:references = "http://ukclimateprojections.metoffice.gov.uk/" ;
		:resolution = "river" ;
		:scenario = "rcp85" ;
		:source = "Probabilistic climate prediction based on family of Met Office Hadley Centre climate models HadCM3, HadRM3 and HadSM3, plus climate models from other climate centres contributing to IPCC AR5 and CFMIP." ;
		:time_slice_type = "1y" ;
		:title = "UKCP18 probabilistic projections for specific humidity anomaly at 1.5m (%) for UK land points, for the RCP 8.5 scenario with a 1981-2000 baseline." ;
		:version = "v20181220" ;
		:Conventions = "CF-1.5" ;
}
