netcdf ESACCI-GHG-L2-CH4-CO-TROPOMI-WFMD-20171110-fv2 {
dimensions:
	sounding_dim = 11254 ;
	level_dim = 21 ;
	layer_dim = 20 ;
	corners_dim = 4 ;
variables:
	double time(sounding_dim) ;
		time:standard_name = "time" ;
		time:long_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00" ;
		time:calendar = "standard" ;
	float latitude(sounding_dim) ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
		latitude:units = "degree_north" ;
		latitude:valid_range = -90.f, 90.f ;
		latitude:comment = "Center latitude of the measurement" ;
	float longitude(sounding_dim) ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
		longitude:units = "degree_east" ;
		longitude:valid_range = -180.f, 180.f ;
		longitude:comment = "Center longitude of the measurement" ;
	float solar_zenith_angle(sounding_dim) ;
		solar_zenith_angle:standard_name = "solar_zenith_angle" ;
		solar_zenith_angle:long_name = "solar_zenith_angle" ;
		solar_zenith_angle:units = "degree" ;
		solar_zenith_angle:comment = "Solar zenith angle is the the angle between the line of sight to the sun and the local vertical." ;
	float sensor_zenith_angle(sounding_dim) ;
		sensor_zenith_angle:standard_name = "sensor_zenith_angle" ;
		sensor_zenith_angle:long_name = "sensor_zenith_angle" ;
		sensor_zenith_angle:units = "degree" ;
		sensor_zenith_angle:comment = "Sensor zenith angle is the the angle between the line of sight to the sensor and the local vertical." ;
	float azimuth_difference(sounding_dim) ;
		azimuth_difference:long_name = "azimuth difference" ;
		azimuth_difference:units = "degree" ;
		azimuth_difference:comment = "Relative azimuth angle between sun and sensor direction." ;
	float xch4(sounding_dim) ;
		xch4:standard_name = "dry_atmosphere_mole_fraction_of_methane" ;
		xch4:long_name = "column-averaged dry air mole fraction of atmospheric methane" ;
		xch4:units = "1e-9" ;
		xch4:comment = "Retrieved column-averaged dry air mole fraction of atmospheric methane (XCH4) in ppb" ;
	float xch4_uncertainty(sounding_dim) ;
		xch4_uncertainty:long_name = "1-sigma uncertainty of the retrieved column-averaged dry air mole fraction of atmospheric methane" ;
		xch4_uncertainty:units = "1e-9" ;
		xch4_uncertainty:comment = "1-sigma uncertainty of the retrieved column-averaged dry air mole fraction of atmospheric methane (XCH4) in ppb" ;
	int xch4_quality_flag(sounding_dim) ;
		xch4_quality_flag:long_name = "quality flag for the retrieved column-averaged dry air mole fraction of atmospheric methane" ;
		xch4_quality_flag:flag_values = 0, 1 ;
		xch4_quality_flag:flag_meanings = "good_quality potentially_bad_quality" ;
		xch4_quality_flag:comment = "0=good, 1=bad" ;
	float xco(sounding_dim) ;
		xco:long_name = "column-averaged dry air mole fraction of atmospheric carbon monoxide" ;
		xco:units = "1e-9" ;
		xco:comment = "Retrieved column-averaged dry air mole fraction of atmospheric carbon monoxide (XCO) in ppb" ;
	float xco_uncertainty(sounding_dim) ;
		xco_uncertainty:long_name = "1-sigma uncertainty of the retrieved column-averaged dry air mole fraction of atmospheric carbon monoxide" ;
		xco_uncertainty:units = "1e-9" ;
		xco_uncertainty:comment = "1-sigma uncertainty of the retrieved column-averaged dry air mole fraction of atmospheric carbon monoxide (XCO) in ppb" ;
	int xco_quality_flag(sounding_dim) ;
		xco_quality_flag:long_name = "quality flag for the retrieved column-averaged dry air mole fraction of atmospheric carbon monoxide" ;
		xco_quality_flag:flag_values = 0, 1 ;
		xco_quality_flag:flag_meanings = "good_quality potentially_bad_quality" ;
		xco_quality_flag:comment = "0=good, 1=bad" ;
	float pressure_levels(sounding_dim, level_dim) ;
		pressure_levels:long_name = "pressure levels" ;
		pressure_levels:units = "hPa" ;
		pressure_levels:comment = "Pressure levels define the boundaries of the averaging kernel and a priori profile layers.\n",
			"Levels are ordered from surface to top of atmosphere." ;
	float pressure_weight(sounding_dim, layer_dim) ;
		pressure_weight:long_name = "pressure weight" ;
		pressure_weight:units = "1" ;
		pressure_weight:comment = "Layer dependent weights needed to apply the averaging kernels." ;
	float ch4_profile_apriori(sounding_dim, layer_dim) ;
		ch4_profile_apriori:long_name = "a priori dry air mole fraction profile of atmospheric methane" ;
		ch4_profile_apriori:units = "1e-9" ;
		ch4_profile_apriori:comment = "A priori dry-air mole fraction profile of atmospheric methane in ppb.\n",
			"All values represent layer averages within the corresponding pressure levels.\n",
			"Profiles are ordered from surface to top of atmosphere." ;
	float xch4_averaging_kernel(sounding_dim, layer_dim) ;
		xch4_averaging_kernel:long_name = "xch4 averaging kernel" ;
		xch4_averaging_kernel:units = "1" ;
		xch4_averaging_kernel:comment = "Represents the altitude sensitivity of the retrieval as a function of pressure.\n",
			"All values represent layer averages within the corresponding pressure levels.\n",
			"Profiles are ordered from surface to top of atmosphere." ;
	float co_profile_apriori(sounding_dim, layer_dim) ;
		co_profile_apriori:long_name = "a priori dry air mole fraction profile of atmospheric carbon monoxide" ;
		co_profile_apriori:units = "1e-9" ;
		co_profile_apriori:comment = "A priori dry-air mole fraction profile of atmospheric carbon monoxide in ppb.\n",
			"All values represent layer averages within the corresponding pressure levels.\n",
			"Profiles are ordered from surface to top of atmosphere." ;
	float xco_averaging_kernel(sounding_dim, layer_dim) ;
		xco_averaging_kernel:long_name = "xco averaging kernel" ;
		xco_averaging_kernel:units = "1" ;
		xco_averaging_kernel:comment = "Represents the altitude sensitivity of the retrieval as a function of pressure.\n",
			"All values represent layer averages within the corresponding pressure levels.\n",
			"Profiles are ordered from surface to top of atmosphere." ;
	int orbit_number(sounding_dim) ;
		orbit_number:long_name = "orbit number" ;
		orbit_number:units = "1" ;
		orbit_number:comment = "Orbit number" ;
	int scanline(sounding_dim) ;
		scanline:long_name = "along track dimension index" ;
		scanline:units = "1" ;
		scanline:comment = "This dimension variable defines the indices along track" ;
	int ground_pixel(sounding_dim) ;
		ground_pixel:long_name = "across track dimension index" ;
		ground_pixel:units = "1" ;
		ground_pixel:comment = "This dimension variable defines the indices across track" ;
	float latitude_corners(sounding_dim, corners_dim) ;
		latitude_corners:long_name = "latitude_corners" ;
		latitude_corners:units = "degree_north" ;
		latitude_corners:valid_range = -90.f, 90.f ;
		latitude_corners:comment = "Corner latitudes of the measurement" ;
	float longitude_corners(sounding_dim, corners_dim) ;
		longitude_corners:long_name = "longitude_corners" ;
		longitude_corners:units = "degree_east" ;
		longitude_corners:valid_range = -180.f, 180.f ;
		longitude_corners:comment = "Corner longitudes of the measurement" ;
	float altitude(sounding_dim) ;
		altitude:standard_name = "altitude" ;
		altitude:long_name = "altitude" ;
		altitude:units = "m" ;
		altitude:comment = "Average surface altitude" ;
	float surface_roughness(sounding_dim) ;
		surface_roughness:long_name = "surface roughness" ;
		surface_roughness:units = "m" ;
		surface_roughness:comment = "Surface roughness" ;
	float apparent_albedo(sounding_dim) ;
		apparent_albedo:long_name = "apparent surface albedo" ;
		apparent_albedo:units = "1" ;
		apparent_albedo:comment = "Retrieved surface albedo at 2313nm" ;
	int land_fraction(sounding_dim) ;
		land_fraction:long_name = "land fraction" ;
		land_fraction:units = "1e-2" ;
		land_fraction:valid_range = 0, 100 ;
		land_fraction:comment = "Land fraction of the observed scene in percent" ;
	float cloud_parameter(sounding_dim) ;
		cloud_parameter:long_name = "cloud parameter from strong water vapour absorption" ;
		cloud_parameter:units = "1" ;
		cloud_parameter:comment = "Ratio of measured to cloud-free reference radiance for selected strong water vapour lines" ;
	float co_column(sounding_dim) ;
		co_column:long_name = "vertical column of carbon monoxide" ;
		co_column:units = "mol m-2" ;
		co_column:multiplication_factor_to_convert_to_molecules_percm2 = 6.022141e+19 ;
		co_column:comment = "Retrieved vertical column amount of carbon monoxide" ;
	float h2o_column(sounding_dim) ;
		h2o_column:long_name = "vertical column of water vapour" ;
		h2o_column:units = "g cm-2" ;
		h2o_column:comment = "Retrieved vertical column amount of water vapour" ;
	float h2o_column_uncertainty(sounding_dim) ;
		h2o_column_uncertainty:long_name = "1-sigma uncertainty of the retrieved vertical column of atmospheric water vapour" ;
		h2o_column_uncertainty:units = "g cm-2" ;
		h2o_column_uncertainty:comment = "1-sigma uncertainty of the retrieved vertical column of atmospheric water vapour" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1.1|hdf5libversion=1.8.18" ;
		:title = "TROPOMI/WFMD XCH4 and XCO" ;
		:institution = "University of Bremen" ;
		:source = "TROPOMI L1B version 01.00.00" ;
		:history = "2021 - product generated with WFMD" ;
		:tracking_id = "6c455a82-fd17-4eee-8e00-46d9ed36a40f" ;
		:Conventions = "CF-1.6" ;
		:product_version = "v1.5" ;
		:summary = "Weighting Function Modified DOAS (WFMD) was adjusted to simultaneously retrieve column-averaged dry air\n",
			"mole fractions of atmospheric methane and carbon monoxide from the shortwave-infrared (SWIR) nadir spectra\n",
			"of the TROPOMI instrument onboard Sentinel-5 Precursor." ;
		:keywords = "satellite, Sentinel-5 Precursor, TROPOMI, atmosphere, methane, carbon monoxide" ;
		:id = "ESACCI-GHG-L2-CH4-CO-TROPOMI-WFMD-20171110-fv2.nc" ;
		:naming_authority = "iup.uni-bremen.de" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD)" ;
		:cdm_data_type = "point" ;
		:comment = "These data were produced at the University of Bremen in the framework of the ESA GHG-CCI project" ;
		:date_created = "20210713T015023Z" ;
		:creator_name = "University of Bremen, IUP, Oliver Schneising" ;
		:creator_email = "schneising@iup.physik.uni-bremen.de" ;
		:project = "Climate Change Initiative - European Space Agency" ;
		:geospatial_lat_min = -90 ;
		:geospatial_lat_max = 90 ;
		:geospatial_lat_units = "degree_north" ;
		:geospatial_lon_min = -180 ;
		:geospatial_lon_max = 180 ;
		:geospatial_lon_units = "degree_east" ;
		:geospatial_vertical_min = 0 ;
		:geospatial_vertical_max = 100000 ;
		:time_coverage_start = "20171110T000000Z" ;
		:time_coverage_end = "20171110T235959Z" ;
		:time_coverage_duration = "P1D" ;
		:time_coverage_resolution = "P1D" ;
		:standard_name_vocabulary = "NetCDF Climate and Forecast (CF) Metadata Conventions Version 1.6" ;
		:license = "ESA CCI Data Policy: free and open access" ;
		:platform = "Sentinel-5 Precursor" ;
		:sensor = "TROPOMI" ;
		:spatial_resolution = "7km x 7km at nadir (typically)" ;
}
