netcdf prsn_rcp85_land-rcm_uk_river_01_ann_198012-208011 {
dimensions:
	ensemble_member = 1 ;
	time = 100 ;
	region = 23 ;
	bnds = 2 ;
	string24 = 24 ;
	string27 = 27 ;
variables:
	float prsn(ensemble_member, time, region) ;
		prsn:standard_name = "snowfall_flux" ;
		prsn:long_name = "Snowfall Flux " ;
		prsn:units = "mm/day" ;
		prsn:description = "Snowfall flux at surface" ;
		prsn:label_units = "mm/day" ;
		prsn:plot_label = "Snowfall flux" ;
		prsn:cell_methods = "time: mean" ;
		prsn:coordinates = "ensemble_member_id geo_region year" ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	char geo_region(region, string24) ;
		geo_region:units = "1" ;
		geo_region:long_name = "River" ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:collection = "land-rcm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2019-09-30T00:00:00" ;
		:domain = "uk" ;
		:frequency = "ann" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "river" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 regional realisation from a set of 12 limited-area Met Office Unified Model Global Atmosphere GA7 models at 12km resolution driven by perturbed variants of the global HadGEM3-GC3.05" ;
		:title = "UKCP18 land projections - 12km regional climate model, snowfall flux over the UK for the RCP 8.5 scenario" ;
		:version = "v20190930" ;
		:Conventions = "CF-1.5" ;
}
