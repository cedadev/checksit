netcdf wsgmax10m_rcp85_land-cpm_uk_2.2km_01_1hr_19801201-19801230 {
dimensions:
	ensemble_member = 1 ;
	time = 720 ;
	grid_latitude = 606 ;
	grid_longitude = 484 ;
	bnds = 2 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float wsgmax10m(ensemble_member, time, grid_latitude, grid_longitude) ;
		wsgmax10m:_FillValue = 1.e+20f ;
		wsgmax10m:standard_name = "wind_speed_of_gust" ;
		wsgmax10m:long_name = "Maximum Wind Speed of Gust at 10m" ;
		wsgmax10m:units = "m s-1" ;
		wsgmax10m:description = "Wind speed gust maximum at 10m" ;
		wsgmax10m:label_units = "m s-1" ;
		wsgmax10m:plot_label = "Wind speed gust maximum (m s-1)" ;
		wsgmax10m:cell_methods = "time: mean" ;
		wsgmax10m:grid_mapping = "rotated_latitude_longitude" ;
		wsgmax10m:coordinates = "ensemble_member_id latitude longitude month_number year yyyymmddhh" ;
	int rotated_latitude_longitude ;
		rotated_latitude_longitude:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_latitude_longitude:longitude_of_prime_meridian = 0. ;
		rotated_latitude_longitude:earth_radius = 6371229. ;
		rotated_latitude_longitude:grid_north_pole_latitude = 37.5 ;
		rotated_latitude_longitude:grid_north_pole_longitude = 177.5 ;
		rotated_latitude_longitude:north_pole_grid_longitude = 0. ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	double grid_latitude(grid_latitude) ;
		grid_latitude:axis = "Y" ;
		grid_latitude:bounds = "grid_latitude_bnds" ;
		grid_latitude:units = "degrees" ;
		grid_latitude:standard_name = "grid_latitude" ;
	double grid_latitude_bnds(grid_latitude, bnds) ;
	double grid_longitude(grid_longitude) ;
		grid_longitude:axis = "X" ;
		grid_longitude:bounds = "grid_longitude_bnds" ;
		grid_longitude:units = "degrees" ;
		grid_longitude:standard_name = "grid_longitude" ;
	double grid_longitude_bnds(grid_longitude, bnds) ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	double latitude(grid_latitude, grid_longitude) ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	double longitude(grid_latitude, grid_longitude) ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;
	char yyyymmddhh(time, string64) ;
		yyyymmddhh:units = "1" ;
		yyyymmddhh:long_name = "yyyymmddhh" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.6.1|hdf5libversion=1.10.4" ;
		:collection = "land-cpm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2021-05-12T10:33:17" ;
		:domain = "uk" ;
		:frequency = "1hr" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "2.2km" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 realisation from a set of 12 convection-permitting models (HadREM3-RA11M) driven by perturbed variants of the Met Office Unified Model Global Atmosphere GA7 model (HadREM3-GA705) at 12km resolution.  The HadREM3-GA705 models were driven by perturbed variants of the global HadGEM3-GC3.05" ;
		:title = "UKCP18 land projections - 2.2km convection-permitting climate model, Maximum Wind Speed of Gust at 10m over the UK for the RCP8.5 scenario" ;
		:version = "v20210615" ;
		:Conventions = "CF-1.7" ;
}
