netcdf sfcWind_rcp85_land-gcm_uk_region_01_day_18991201-20991130 {
dimensions:
	ensemble_member = 1 ;
	time = 72000 ;
	region = 16 ;
	bnds = 2 ;
	string24 = 24 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float sfcWind(ensemble_member, time, region) ;
		sfcWind:standard_name = "wind_speed" ;
		sfcWind:long_name = "Wind speed at 10m" ;
		sfcWind:units = "m s-1" ;
		sfcWind:description = "Wind speed" ;
		sfcWind:label_units = "m s-1" ;
		sfcWind:plot_label = "Wind speed at 10m (m s-1)" ;
		sfcWind:cell_methods = "time: mean" ;
		sfcWind:coordinates = "ensemble_member_id geo_region month_number year yyyymmdd" ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	char geo_region(region, string24) ;
		geo_region:units = "1" ;
		geo_region:long_name = "Region" ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;
	char yyyymmdd(time, string64) ;
		yyyymmdd:units = "1" ;
		yyyymmdd:long_name = "yyyymmdd" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.4.1|hdf5libversion=1.8.17" ;
		:collection = "land-gcm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2018-11-10T15:52:53" ;
		:domain = "uk" ;
		:frequency = "day" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "region" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 global realisation from a set of 15 perturbed variants of HadGEM3-GC3.05 and 13 CMIP5 members that passed a qualitative evaluation" ;
		:title = "UKCP18 land projections - 60km global climate model, wind speed at 10m (m s-1) over the UK for the RCP 8.5 scenario" ;
		:version = "v20181122" ;
		:Conventions = "CF-1.5" ;
}
