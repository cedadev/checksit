netcdf pr_rcp85_land-cpm_uk_river_01_seas-20y_198012-200011 {
dimensions:
	ensemble_member = 1 ;
	time = 4 ;
	region = 23 ;
	bnds = 2 ;
	string21 = 21 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float pr(ensemble_member, time, region) ;
		pr:_FillValue = 1.e+20f ;
		pr:standard_name = "lwe_precipitation_rate" ;
		pr:long_name = "Precipitation rate" ;
		pr:units = "mm/day" ;
		pr:description = "Precipitation rate" ;
		pr:label_units = "mm/day" ;
		pr:plot_label = "Precipitation rate (mm/day)" ;
		pr:cell_methods = "time: mean" ;
		pr:coordinates = "ensemble_member_id geo_region season year" ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	char geo_region(region, string21) ;
		geo_region:units = "1" ;
		geo_region:long_name = "River" ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	char season(time, string64) ;
		season:units = "1" ;
		season:long_name = "season" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:_NCProperties = "version=2,netcdf=4.6.3,hdf5=1.10.5" ;
		:collection = "land-cpm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2021-06-15T00:00:00" ;
		:domain = "uk" ;
		:frequency = "seas-20y" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "river" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 realisation from a set of 12 convection-permitting models (HadREM3-RA11M) driven by perturbed variants of the Met Office Unified Model Global Atmosphere GA7 model (HadREM3-GA705) at 12km resolution. The HadREM3-GA705 models were driven by perturbed variants of the global HadGEM3-GC3.05" ;
		:title = "UKCP18 land projections - 2.2km convection-permitting climate model regionally-averaged,  precipitation rate (mm/day) over the UK for the RCP 8.5 scenario" ;
		:version = "v20210615" ;
		:Conventions = "CF-1.7" ;
}
