netcdf clt_rcp85_land-cpm_uk_5km_01_ann-20y_198012-199011 {

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.6.1|hdf5libversion=1.10.4" ;
}
