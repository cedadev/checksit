netcdf tasAnom_rcp85_land-prob_uk_country_sample_b8100_1y_seas_19601201-20991130 {
dimensions:
	time = UNLIMITED ; // (556 currently)
	region = 8 ;
	sample = 3000 ;
	bnds = 2 ;
	string24 = 24 ;
	string64 = 64 ;
variables:
	float tasAnom(time, region, sample) ;
		tasAnom:standard_name = "air_temperature" ;
		tasAnom:long_name = "Mean air temperature" ;
		tasAnom:units = "degC" ;
		tasAnom:anomaly_type = "absolute_change" ;
		tasAnom:description = "Mean air temperature" ;
		tasAnom:label_units = "°C" ;
		tasAnom:plot_label = "Mean air temperature anomaly at 1.5m (°C)" ;
		tasAnom:cell_methods = "time: mean" ;
		tasAnom:coordinates = "geo_region season year" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	int sample(sample) ;
		sample:units = "1" ;
		sample:long_name = "sample" ;
	char geo_region(region, string24) ;
		geo_region:units = "1" ;
		geo_region:long_name = "Country" ;
	char season(time, string64) ;
		season:units = "1" ;
		season:long_name = "season" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:baseline_period = "b8100" ;
		:collection = "land-prob" ;
		:contact = "ukcpproject@metoffice.gov.uk, UKCP Team, Met Office Hadley Centre" ;
		:creation_date = "2018-12-23T15:59:37" ;
		:domain = "uk" ;
		:frequency = "seas" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:prob_data_type = "sample" ;
		:project = "UKCP18" ;
		:references = "http://ukclimateprojections.metoffice.gov.uk/" ;
		:resolution = "country" ;
		:scenario = "rcp85" ;
		:source = "Probabilistic climate prediction based on family of Met Office Hadley Centre climate models HadCM3, HadRM3 and HadSM3, plus climate models from other climate centres contributing to IPCC AR5 and CFMIP." ;
		:time_slice_type = "1y" ;
		:title = "UKCP18 probabilistic projections for mean air temperature anomaly at 1.5m (K) for UK land points, for the RCP 8.5 scenario with a 1981-2000 baseline." ;
		:version = "v20181220" ;
		:Conventions = "CF-1.5" ;
}
