netcdf prsn_rcp85_land-cpm_uk_5km_01_seas-20y_198012-200011 {
dimensions:
	ensemble_member = 1 ;
	time = 4 ;
	projection_y_coordinate = 244 ;
	projection_x_coordinate = 180 ;
	bnds = 2 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float prsn(ensemble_member, time, projection_y_coordinate, projection_x_coordinate) ;
		prsn:_FillValue = 1.e+20f ;
		prsn:standard_name = "snowfall_flux" ;
		prsn:long_name = "Snowfall Flux " ;
		prsn:units = "mm/day" ;
		prsn:description = "Snowfall flux at surface" ;
		prsn:label_units = "mm/day" ;
		prsn:plot_label = "Snowfall flux" ;
		prsn:cell_methods = "time: mean" ;
		prsn:grid_mapping = "transverse_mercator" ;
		prsn:coordinates = "ensemble_member_id latitude longitude season year" ;
	int transverse_mercator ;
		transverse_mercator:grid_mapping_name = "transverse_mercator" ;
		transverse_mercator:longitude_of_prime_meridian = 0. ;
		transverse_mercator:semi_major_axis = 6377563.396 ;
		transverse_mercator:semi_minor_axis = 6356256.909 ;
		transverse_mercator:longitude_of_central_meridian = -2. ;
		transverse_mercator:latitude_of_projection_origin = 49. ;
		transverse_mercator:false_easting = 400000. ;
		transverse_mercator:false_northing = -100000. ;
		transverse_mercator:scale_factor_at_central_meridian = 0.9996012717 ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	double projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:axis = "Y" ;
		projection_y_coordinate:bounds = "projection_y_coordinate_bnds" ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
	double projection_y_coordinate_bnds(projection_y_coordinate, bnds) ;
	double projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:axis = "X" ;
		projection_x_coordinate:bounds = "projection_x_coordinate_bnds" ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
	double projection_x_coordinate_bnds(projection_x_coordinate, bnds) ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	double latitude(projection_y_coordinate, projection_x_coordinate) ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
	double longitude(projection_y_coordinate, projection_x_coordinate) ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
	char season(time, string64) ;
		season:units = "1" ;
		season:long_name = "season" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:_NCProperties = "version=2,netcdf=4.6.3,hdf5=1.10.5" ;
		:collection = "land-cpm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2021-06-15T00:00:00" ;
		:domain = "uk" ;
		:frequency = "seas-20y" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "5km" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 realisation from a set of 12 convection-permitting models (HadREM3-RA11M) driven by perturbed variants of the Met Office Unified Model Global Atmosphere GA7 model (HadREM3-GA705) at 12km resolution. The HadREM3-GA705 models were driven by perturbed variants of the global HadGEM3-GC3.05" ;
		:title = "UKCP18 land projections - 2.2km convection-permitting climate model regridded to 5km, snowfall flux over the UK for the RCP 8.5 scenario" ;
		:version = "v20210615" ;
		:Conventions = "CF-1.7" ;
}
