netcdf ESACCI-GHG-L2-CO2-GOSAT2-SRFP-20191231-fv2 {
dimensions:
	sounding_dim = 3393 ;
	polarization_dim = 2 ;
	level_dim = 13 ;
	layer_dim = 12 ;
	window_dim = 4 ;
	char_l1bname = 28 ;
	gain_dim = 6 ;
variables:
	float solar_zenith_angle(sounding_dim) ;
		solar_zenith_angle:long_name = "solar zenith angle" ;
		solar_zenith_angle:units = "degrees" ;
		solar_zenith_angle:comment = "Solar zenith angle is the angle between the line of sight to the sun and the local vertical." ;
	float sensor_zenith_angle(sounding_dim) ;
		sensor_zenith_angle:long_name = "sensor zenith angle" ;
		sensor_zenith_angle:units = "degrees" ;
		sensor_zenith_angle:comment = "Sensor zenith angle is the angle between the line of sight to the sensor and the local vertical." ;
	double time(sounding_dim) ;
		time:long_name = "time" ;
		time:units = "seconds since 1970-01-01 00:00:00" ;
		time:calender = "standard" ;
	float longitude(sounding_dim) ;
		longitude:long_name = "longitude" ;
		longitude:units = "degrees_east" ;
		longitude:comment = "Center longitude of the measurement." ;
		longitude:valid_range = -180., 180. ;
	float latitude(sounding_dim) ;
		latitude:long_name = "latitude" ;
		latitude:units = "degrees_north" ;
		latitude:comment = "Center latitude of the measurement." ;
		latitude:valid_range = -90., 90. ;
	float pressure_levels(sounding_dim, level_dim) ;
		pressure_levels:long_name = "pressure_levels" ;
		pressure_levels:units = "hPa" ;
		pressure_levels:comment = "Pressure levels define the boundaries of the averaging kernel and mole fraction profile layers. Surface pressure is represented by the 1st element, i.e., profiles are ordered from surface to top of atmosphere." ;
	float pressure_weight(sounding_dim, layer_dim) ;
		pressure_weight:long_name = "pressure weight" ;
		pressure_weight:units = "1" ;
		pressure_weight:comment = "Pressure weights are the layer dependent weights needed to apply the averaging kernels." ;
	float xco2(sounding_dim) ;
		xco2:long_name = "column-average dry-air mole fraction of atmospheric carbon dioxide" ;
		xco2:units = "1e-9" ;
		xco2:comment = "Retrieved column-average dry-air mole fraction of atmospheric carbon dioxide (XCO2) in ppm." ;
	float xco2_uncertainty(sounding_dim) ;
		xco2_uncertainty:long_name = "1-sigma uncertainty of the retrieved column-average dry-air mole fraction of atmospheric carbon dioxide" ;
		xco2_uncertainty:units = "1e-9" ;
		xco2_uncertainty:comment = "1-sigma uncertainty of the retrieved column-average dry-air mole fraction of atmospheric carbon dioxide (XCO2) in ppm." ;
	float xco2_averaging_kernel(sounding_dim, layer_dim) ;
		xco2_averaging_kernel:long_name = "normalized column averaging kernel" ;
		xco2_averaging_kernel:units = "1" ;
		xco2_averaging_kernel:comment = "The normalized column-averaging kernel represents the sensitivity of the retrieved XCO2 to the atmospheric carbon dioxide mole fraction depending on pressure (height). All values represent layer averages within the corresponding pressure levels. Values near one are ideal and indicate that the influence of the a priori is minimal. Profiles are ordered from surface to top of atmosphere." ;
	float co2_profile_apriori(sounding_dim, layer_dim) ;
		co2_profile_apriori:long_name = "a priori dry-air mole fraction profile of atmospheric carbon dioxide" ;
		co2_profile_apriori:units = "1e-9" ;
		co2_profile_apriori:comment = "A priori dry-air mole fraction profile of atmospheric carbon dioxide in ppm (http://www.atmos-meas-tech.net/5/1349/2012/amt-5-1349-2012.html). All values represent layer averages within the corresponding pressure levels. Profiles are ordered from surface to top of atmosphere." ;
	int xco2_quality_flag(sounding_dim) ;
		xco2_quality_flag:long_name = "xco2_quality flag" ;
		xco2_quality_flag:units = "1" ;
		xco2_quality_flag:values = "0B, 1B; // byte" ;
		xco2_quality_flag:meanings = "Quality flag for XCO2 retrieval" ;
		xco2_quality_flag:comment = "0=good, 1=bad" ;
	int flag_landtype(sounding_dim) ;
		flag_landtype:long_name = "flag for land / ocean soundings" ;
		flag_landtype:units = "1" ;
		flag_landtype:comment = "0 = no glint, 1 = glint" ;
	int flag_sunglint(sounding_dim) ;
		flag_sunglint:long_name = "flag for normal / sunglint soundings" ;
		flag_sunglint:units = "1" ;
		flag_sunglint:comment = "0 = no glint, 1 = glint" ;
	char gain(sounding_dim, gain_dim) ;
		gain:long_name = "gain" ;
		gain:units = "1" ;
		gain:comment = "Number of gain coefficient is stored for each band. The gain coefficient of each band is calculated from solar calibration mode data. The order is 1P, 1S, 2P, 2S, 3P, 3S." ;
	int exposure_id(sounding_dim) ;
		exposure_id:long_name = "exposure id" ;
		exposure_id:units = "1" ;
		exposure_id:comment = "Exposure identification number of the sounding" ;
	char l1b_name(sounding_dim, char_l1bname) ;
		l1b_name:long_name = "level 1B name" ;
		l1b_name:units = "1" ;
		l1b_name:comment = "Name of the Level 1B file of the sounding" ;
	float signal_to_noise_window(sounding_dim, polarization_dim, window_dim) ;
		signal_to_noise_window:long_name = "signal to noise ratio" ;
		signal_to_noise_window:units = "1" ;
		signal_to_noise_window:comment = "The signal to noise ratio per retrieval window for both polarization directions. Window 1 ranges between 757 nm and 773 nm, Window 2 ranges between 1.59 um and 1.62 um, Window 3 ranges between 1.63 um and 1.65 um and Window 4 ranges between 2.04 um and 2.08 um" ;
	float dry_airmass_layer(sounding_dim, layer_dim) ;
		dry_airmass_layer:long_name = "Dry airmass per layer" ;
		dry_airmass_layer:units = "m-2" ;
		dry_airmass_layer:comment = "The dry airmass per layer, units are molecules m-2" ;
	float altitude(sounding_dim) ;
		altitude:long_name = "Altitude" ;
		altitude:units = "m" ;
		altitude:comment = "Altitude is the surface elevation in meters" ;
	float air_temperature(sounding_dim, level_dim) ;
		air_temperature:long_name = "Air temperature at each level" ;
		air_temperature:units = "K" ;
		air_temperature:comment = "" ;
	float surface_altitude_stdv(sounding_dim) ;
		surface_altitude_stdv:long_name = "Standard deviation of the surface elevation" ;
		surface_altitude_stdv:units = "m" ;
		surface_altitude_stdv:comment = "Standard deviation of the surface elevation within the area of the GOSAT-2 sounding, as derived from the SRTM database" ;
	float x_wind(sounding_dim, level_dim) ;
		x_wind:long_name = "grid_eastward_wind " ;
		x_wind:units = "m s-1" ;
		x_wind:comment = "\'x\' indicates a vector component along the grid x-axis, positive with increasing x. Wind is defined as a two-dimensional (horizontal) air velocity vector, with no vertical component. (Vertical motion in the atmosphere has the standard name upward_air_velocity.)" ;
	float y_wind(sounding_dim, level_dim) ;
		y_wind:long_name = "grid_northward_wind" ;
		y_wind:units = "m s-1" ;
		y_wind:comment = "\'y\' indicates a vector component along the grid y-axis, positive with increasing y. Wind is defined as a two-dimensional (horizontal) air velocity vector, with no vertical component. (Vertical motion in the atmosphere has the standard name upward_air_velocity.) " ;
	float chi2(sounding_dim) ;
		chi2:long_name = "Chi-squared" ;
		chi2:unit = "1" ;
		chi2:comment = "Chi_squared value of the sounding" ;
	float optical_thickness_of_atmosphere_layer_due_to_ambient_aerosol(sounding_dim, window_dim) ;
		optical_thickness_of_atmosphere_layer_due_to_ambient_aerosol:long_name = "Aerosol optical thickness per retrieval window" ;
		optical_thickness_of_atmosphere_layer_due_to_ambient_aerosol:unit = "1" ;
		optical_thickness_of_atmosphere_layer_due_to_ambient_aerosol:comment = "\'Layer\' means any layer with upper and lower boundaries that have constant values in some vertical coordinate. There must be a vertical coordinate variable indicating the extent of the layer(s). If the layers are model layers, the vertical coordinate can be model_level_number, but it is recommended to specify a physical coordinate (in a scalar or auxiliary coordinate variable) as well. The optical thickness is the integral along the path of radiation of a volume scattering/absorption/attenuation coefficient. The radiative flux is reduced by a factor exp(-optical_thickness) on traversing the path. A coordinate variable of radiation_wavelength or radiation_frequency can be specified to indicate that the optical thickness applies at specific wavelengths or frequencies. \'Aerosol\' means the suspended liquid or solid particles in air (except cloud droplets). \'Ambient aerosol\' is aerosol that has taken up ambient water through hygroscopic growth. The extent of hygroscopic growth depends on the relative humidity and the composition of the aerosol. The specification of a physical process by the phrase due_to_process means that the quantity named is a single term in a sum of terms which together compose the general quantity named by omitting the phrase. Window 1 ranges between 757 nm and 773 nm, window 2 ranges from 1.59 um and 1.62 um, window 3 ranges between 1.63 um and 1.65 um and window 4 ranges between 2.04 um and 2.08 um" ;
	float raw_xco2(sounding_dim) ;
		raw_xco2:long_name = "Raw retrieved XCO2 column" ;
		raw_xco2:units = "1e-9" ;
		raw_xco2:comment = "The retrieved raw XCO2 total column before bias correction" ;
	float raw_xco2_err(sounding_dim) ;
		raw_xco2_err:long_name = "Raw uncertainty on the XCO2 total column" ;
		raw_xco2_err:units = "1e-9" ;
		raw_xco2_err:commment = "The raw uncertainty due to measurement noise on the XCO2 total column" ;
	float h2o_column(sounding_dim) ;
		h2o_column:long_name = "H2O total column" ;
		h2o_column:units = "m-2" ;
		h2o_column:comment = "The retrieved H2O total column in units of molecules m-2" ;
	float surface_albedo_758(sounding_dim) ;
		surface_albedo_758:long_name = "Surface albedo at 758 nm" ;
		surface_albedo_758:units = "1" ;
		surface_albedo_758:comment = "The retrieved surface albedo for window 1, at 758 nm" ;
	float surface_albedo_1593(sounding_dim) ;
		surface_albedo_1593:long_name = "Surface albedo at 1593 nm" ;
		surface_albedo_1593:units = "1" ;
		surface_albedo_1593:comment = "The retrieved surface albedo for window 2, at 1593 nm" ;
	float surface_albedo_1629(sounding_dim) ;
		surface_albedo_1629:long_name = "Surface albedo at 1629 nm" ;
		surface_albedo_1629:units = "1" ;
		surface_albedo_1629:comment = "The retrieved surface albedo for window 3, at 1629 nm" ;
	float surface_albedo_2042(sounding_dim) ;
		surface_albedo_2042:long_name = "Surface albedo at 2042 nm" ;
		surface_albedo_2042:units = "1" ;
		surface_albedo_2042:comment = "The retrieved surface albedo for window 4, at 2042 nm" ;
	float intensity_offset_o2a(sounding_dim) ;
		intensity_offset_o2a:long_name = "Intensity offset in the O2A-band" ;
		intensity_offset_o2a:units = "W cm-2" ;
		intensity_offset_o2a:comment = "The retrieved intensity offset in the O2A-band" ;
	float aerosol_size(sounding_dim) ;
		aerosol_size:long_name = "Retrieved size parameter of the aerosol distribution" ;
		aerosol_size:units = "1" ;
		aerosol_size:comment = "The size parameter is the exponent of the power-law slope of the aerosol size distribution" ;
	float aerosol_central_height(sounding_dim) ;
		aerosol_central_height:long_name = "Retrieved aerosol peak height" ;
		aerosol_central_height:units = "m" ;
		aerosol_central_height:comment = "Peak height of the aerosol Gaussian height distribution" ;
	float aerosol_total_column(sounding_dim) ;
		aerosol_total_column:long_name = "Retrieved aerosol total column" ;
		aerosol_total_column:units = "m-2" ;
		aerosol_total_column:comment = "The retrieved total aerosol column in units of particles m-2" ;

// global attributes:
		:title = "ESA CCI GOSAT2 SRFP XCO2" ;
		:institution = "SRON Netherlands Institute for Space Research" ;
		:source = "GOSAT2 L1B version v210" ;
		:history = "02.11.2022 -  product generated with RemoTeC v2.0.0" ;
		:references = "http://www.esa-ghg-cii.org/ \n http://onlinelibrary.wiley.com/doi/10.1002/jgrd.50332/abstract \n http://onlinelibrary.wiley.com/doi/10.1029/2011GL047888/abstract" ;
		:tracking_id = "ea60bd02-6c38-11e5-82fb-d3dc42d9b150" ;
		:Conventions = "CF-1.6" ;
		:product_version = "v2.0.0" ;
		:summary = "The RemoTeC algorithm was designed to analyze GOSAT2 TANSO-FTS2 data, both for CO2 and CH4. It utilizes both a PROXY approach (for CH4) where the scattering due to clouds and aerosols is taken into account by multiplying the observed ratio of CH4/CO2 with a prior model CO2, as well as a Full Physics approach (for CH4 and CO2) where the CO2 and CH4 spectra are simultaneously fitted with aerosol parameters to retrieve the scattering information due to clouds and aerosols. This product uses the Full Physics approach for CH4 " ;
		:keywords = "satellite, GOSAT2, TANSO-FTS2, atmosphere, carbondioxide" ;
		:id = "ESACCI-GHG-L2-CO2-GOSAT2-SRFP-20191231-fv2.nc" ;
		:naming_authority = "home.sron.nl" ;
		:keywords_vocabulary = "NASA Global Change Master Directory (GCMD)" ;
		:cdm_data_type = "point" ;
		:comment = "These data were produced at SRON Netherlands Institute for Space Research in the frame of the ESA GHG CCI project" ;
		:date_created = "CreatedWed Nov  2 09:32:11 2022" ;
		:creator_name = "SRON Netherlands Institute for Space Research, Andrew Barr" ;
		:creator_url = "ftp://ftp.sron.nl/pub/pub/RemoTeC/" ;
		:creator_email = "a.g.barr@sron.nl" ;
		:project = "Climate Change Initiative - European Space Agency" ;
		:geospatial_lat_min = "-90.0f; // float" ;
		:geospatial_lat_max = "90.0f; // float" ;
		:geospatial_lat_units = "degrees_north" ;
		:geospatial_lon_min = "-180.0f; // float" ;
		:geospatial_lon_max = "180.0f; // float" ;
		:geospatial_lon_units = "degrees_east" ;
		:geospatial_vertical_min = "0.0f; // float" ;
		:geospatial_vertical_max = "100000.0; // float" ;
		:time_coverage_start = "20191231T000000Z" ;
		:time_coverage_end = "20191231T235959Z" ;
		:time_coverage_duration = "P1D" ;
		:time_coverage_resolution = "P1D" ;
		:standard_name_vocabulary = "CF Standard Name Table v79" ;
		:license = "ESA CCI Data Policy: free and open access" ;
		:platform = "GOSAT2" ;
		:sensor = "TANSO-FTS2" ;
		:spatial_resolution = "10.5km x 10.5km at nadir (typically)" ;
		:_CoordSysBuilder = "ucar.nc2.dataset.conv.CF1Convention" ;
}
