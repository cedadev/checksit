netcdf beta_rcp85_land-rcm_eur_12km_01_mon_198012-208011 {
dimensions:
	ensemble_member = 1 ;
	time = 1200 ;
	grid_latitude = 406 ;
	grid_longitude = 418 ;
	bnds = 2 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float beta(ensemble_member, time, grid_latitude, grid_longitude) ;
		beta:_FillValue = 1.e+20f ;
		beta:long_name = "Soil moisture stress factor" ;
		beta:units = "1" ;
		beta:cell_methods = "depth: sum" ;
		beta:grid_mapping = "rotated_latitude_longitude" ;
		beta:coordinates = "ensemble_member_id month_number year yyyymm" ;
	int rotated_latitude_longitude ;
		rotated_latitude_longitude:grid_mapping_name = "rotated_latitude_longitude" ;
		rotated_latitude_longitude:longitude_of_prime_meridian = 0. ;
		rotated_latitude_longitude:earth_radius = 6371229. ;
		rotated_latitude_longitude:grid_north_pole_latitude = 39.25 ;
		rotated_latitude_longitude:grid_north_pole_longitude = 198. ;
		rotated_latitude_longitude:north_pole_grid_longitude = 0. ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	double grid_latitude(grid_latitude) ;
		grid_latitude:axis = "Y" ;
		grid_latitude:bounds = "grid_latitude_bnds" ;
		grid_latitude:units = "degrees" ;
		grid_latitude:standard_name = "grid_latitude" ;
	double grid_latitude_bnds(grid_latitude, bnds) ;
	double grid_longitude(grid_longitude) ;
		grid_longitude:axis = "X" ;
		grid_longitude:bounds = "grid_longitude_bnds" ;
		grid_longitude:units = "degrees" ;
		grid_longitude:standard_name = "grid_longitude" ;
	double grid_longitude_bnds(grid_longitude, bnds) ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;
	char yyyymm(time, string64) ;
		yyyymm:units = "1" ;
		yyyymm:long_name = "yyyymm" ;

// global attributes:
		:_NCProperties = "version=2,netcdf=4.6.3,hdf5=1.10.5" ;
		:collection = "land-rcm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2020-05-31T00:00:00" ;
		:description = "Soil moisture stress factor" ;
		:domain = "eur" ;
		:frequency = "mon" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:label_units = "dimensionless" ;
		:plot_label = "Soil moisture stress factor (dimensionless)" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "12km" ;
		:scenario = "rcp85" ;
		:source = "UKCP18 regional realisation from a set of 12 limited-area Met Office Unified Model Global Atmosphere GA7 models at 12km resolution driven by perturbed variants of the global HadGEM3-GC3.05" ;
		:title = "UKCP18 land projections - 12km regional climate model for the RCP 8.5 scenario" ;
		:version = "v20200531" ;
		:Conventions = "CF-1.7" ;
}
