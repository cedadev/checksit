netcdf rlsAnom_rcp85_land-prob_uk_25km_cdf_b6190_30y_mon_20091201-20991130 {
dimensions:
	time = 84 ;
	projection_y_coordinate = 52 ;
	projection_x_coordinate = 39 ;
	percentile = 111 ;
	bnds = 2 ;
	string64 = 64 ;
variables:
	float rlsAnom(time, projection_y_coordinate, projection_x_coordinate, percentile) ;
		rlsAnom:long_name = "Net Surface long wave flux" ;
		rlsAnom:units = "W m-2" ;
		rlsAnom:anomaly_type = "absolute_change" ;
		rlsAnom:description = "Net Surface long wave flux" ;
		rlsAnom:label_units = "W m-2" ;
		rlsAnom:plot_label = "Net Surface long wave flux anomaly (W m-2)" ;
		rlsAnom:cell_methods = "time: mean" ;
		rlsAnom:grid_mapping = "transverse_mercator" ;
		rlsAnom:coordinates = "latitude longitude month_number season season_year year" ;
	int transverse_mercator ;
		transverse_mercator:grid_mapping_name = "transverse_mercator" ;
		transverse_mercator:longitude_of_prime_meridian = 0. ;
		transverse_mercator:semi_major_axis = 6377563.396 ;
		transverse_mercator:semi_minor_axis = 6356256.909 ;
		transverse_mercator:longitude_of_central_meridian = -2. ;
		transverse_mercator:latitude_of_projection_origin = 49. ;
		transverse_mercator:false_easting = 400000. ;
		transverse_mercator:false_northing = -100000. ;
		transverse_mercator:scale_factor_at_central_meridian = 0.9996012717 ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	double projection_y_coordinate(projection_y_coordinate) ;
		projection_y_coordinate:axis = "Y" ;
		projection_y_coordinate:bounds = "projection_y_coordinate_bnds" ;
		projection_y_coordinate:units = "m" ;
		projection_y_coordinate:standard_name = "projection_y_coordinate" ;
	double projection_y_coordinate_bnds(projection_y_coordinate, bnds) ;
	double projection_x_coordinate(projection_x_coordinate) ;
		projection_x_coordinate:axis = "X" ;
		projection_x_coordinate:bounds = "projection_x_coordinate_bnds" ;
		projection_x_coordinate:units = "m" ;
		projection_x_coordinate:standard_name = "projection_x_coordinate" ;
	double projection_x_coordinate_bnds(projection_x_coordinate, bnds) ;
	double percentile(percentile) ;
		percentile:units = "%" ;
		percentile:long_name = "percentile" ;
	double latitude(projection_y_coordinate, projection_x_coordinate) ;
		latitude:units = "degrees_north" ;
		latitude:standard_name = "latitude" ;
		latitude:long_name = "latitude" ;
	double longitude(projection_y_coordinate, projection_x_coordinate) ;
		longitude:units = "degrees_east" ;
		longitude:standard_name = "longitude" ;
		longitude:long_name = "longitude" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	char season(time, string64) ;
		season:units = "1" ;
		season:long_name = "season" ;
	int season_year(time) ;
		season_year:units = "1" ;
		season_year:long_name = "season_year" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:baseline_period = "b6190" ;
		:collection = "land-prob" ;
		:contact = "ukcpproject@metoffice.gov.uk, UKCP Team, Met Office Hadley Centre" ;
		:creation_date = "2018-10-08T08:34:12" ;
		:domain = "uk" ;
		:frequency = "mon" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:prob_data_type = "cdf" ;
		:project = "UKCP18" ;
		:references = "http://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "25km" ;
		:scenario = "rcp85" ;
		:source = "Probabilistic climate prediction based on family of Met Office Hadley Centre climate models HadCM3, HadRM3 and HadSM3, plus climate models from other climate centres contributing to IPCC AR5 and CFMIP." ;
		:time_slice_type = "30y" ;
		:title = "UKCP18 probabilistic projections for net surface long wave flux anomaly (W m-2) for UK land points, for the RCP 8.5 scenario with a 1961-1990 baseline." ;
		:version = "v20181122" ;
		:Conventions = "CF-1.5" ;
}
