netcdf tasminAnom_rcp85_land-prob_uk_region_pdf_b8100_1y_ann_19601201-20991130 {
dimensions:
	time = UNLIMITED ; // (139 currently)
	region = 16 ;
	percentile = 111 ;
	bnds = 2 ;
	string26 = 26 ;
variables:
	float tasminAnom(time, region, percentile) ;
		tasminAnom:long_name = "Minimum air temperature probability density" ;
		tasminAnom:units = "degC-1" ;
		tasminAnom:anomaly_type = "absolute_change" ;
		tasminAnom:description = "Minimum air temperature" ;
		tasminAnom:label_units = "°C-1" ;
		tasminAnom:plot_label = "Probability density for minimum air temperature anomaly at 1.5m (°C-1)" ;
		tasminAnom:cell_methods = "time: mean" ;
		tasminAnom:coordinates = "geo_region year" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	double percentile(percentile) ;
		percentile:units = "%" ;
		percentile:long_name = "percentile" ;
	char geo_region(region, string26) ;
		geo_region:units = "1" ;
		geo_region:long_name = "Administrative Region" ;
	int year(time) ;
		year:units = "1" ;
		year:long_name = "year" ;

// global attributes:
		:baseline_period = "b8100" ;
		:collection = "land-prob" ;
		:contact = "ukcpproject@metoffice.gov.uk, UKCP Team, Met Office Hadley Centre" ;
		:creation_date = "2018-12-23T16:07:17" ;
		:domain = "uk" ;
		:frequency = "ann" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:prob_data_type = "pdf" ;
		:project = "UKCP18" ;
		:references = "http://ukclimateprojections.metoffice.gov.uk/" ;
		:resolution = "region" ;
		:scenario = "rcp85" ;
		:source = "Probabilistic climate prediction based on family of Met Office Hadley Centre climate models HadCM3, HadRM3 and HadSM3, plus climate models from other climate centres contributing to IPCC AR5 and CFMIP." ;
		:time_slice_type = "1y" ;
		:title = "UKCP18 probabilistic projections for minimum air temperature anomaly at 1.5m (K) for UK land points, for the RCP 8.5 scenario with a 1981-2000 baseline." ;
		:version = "v20181220" ;
		:Conventions = "CF-1.5" ;
}
