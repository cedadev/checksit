netcdf evspsbl_rcp26_land-gcm_uk_region_01_mon-30y_196012-199011 {
dimensions:
	ensemble_member = 1 ;
	time = 12 ;
	region = 16 ;
	bnds = 2 ;
	string20 = 20 ;
	string27 = 27 ;
	string64 = 64 ;
variables:
	float evspsbl(ensemble_member, time, region) ;
		evspsbl:standard_name = "water_evaporation_flux" ;
		evspsbl:long_name = "Evaporation rate" ;
		evspsbl:units = "mm/day" ;
		evspsbl:description = "Evaporation rate" ;
		evspsbl:label_units = "mm/day" ;
		evspsbl:plot_label = "Evaporation rate (mm/day)" ;
		evspsbl:cell_methods = "time: mean" ;
		evspsbl:coordinates = "ensemble_member_id geo_region month_number yyyymm" ;
	int ensemble_member(ensemble_member) ;
		ensemble_member:units = "1" ;
		ensemble_member:long_name = "ensemble_member" ;
	double time(time) ;
		time:axis = "T" ;
		time:bounds = "time_bnds" ;
		time:units = "hours since 1970-01-01 00:00:00" ;
		time:standard_name = "time" ;
		time:calendar = "360_day" ;
	double time_bnds(time, bnds) ;
	int region(region) ;
		region:units = "1" ;
		region:standard_name = "region" ;
	char geo_region(region, string20) ;
		geo_region:units = "1" ;
		geo_region:long_name = "Region" ;
	char ensemble_member_id(ensemble_member, string27) ;
		ensemble_member_id:units = "1" ;
		ensemble_member_id:long_name = "ensemble_member_id" ;
	int month_number(time) ;
		month_number:units = "1" ;
		month_number:long_name = "month_number" ;
	char yyyymm(time, string64) ;
		yyyymm:units = "1" ;
		yyyymm:long_name = "yyyymm" ;

// global attributes:
		:_NCProperties = "version=1|netcdflibversion=4.6.1|hdf5libversion=1.10.4" ;
		:collection = "land-gcm" ;
		:contact = "ukcpproject@metoffice.gov.uk" ;
		:creation_date = "2020-03-02T00:00:00" ;
		:domain = "uk" ;
		:frequency = "mon-30y" ;
		:institution = "Met Office Hadley Centre (MOHC), FitzRoy Road, Exeter, Devon, EX1 3PB, UK." ;
		:institution_id = "MOHC" ;
		:project = "UKCP18" ;
		:references = "https://ukclimateprojections.metoffice.gov.uk" ;
		:resolution = "region" ;
		:scenario = "rcp26" ;
		:source = "UKCP18 global realisation from a set of 15 perturbed variants of HadGEM3-GC3.05 and 13 CMIP5 members that passed a qualitative evaluation" ;
		:title = "UKCP18 land projections - 60km global climate model evaporation rate (mm/day) over the UK for the RCP 8.5 scenario" ;
		:version = "v20200302" ;
		:Conventions = "CF-1.5" ;
}
